`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: ITCR 
// Engineer: ADRIAN CERVANTES SEGURA 
// 
// Create Date: 03.03.2016 01:49:40
// Design Name: 
// Module Name: LUT_SHIFT
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module LUT_SHIFT #(parameter P = 32, parameter D = 5) ( 

input wire CLK, 
input wire EN_ROM1,
input wire [D-1:0] ADRS,
output reg [P-1:0] O_D
);
   
always @(posedge CLK)
      if (EN_ROM1)
         case (ADRS)
            5'b00000: O_D <= 32'b00111111011111110000000000000000;//1-2^(-6-2)
            5'b00001: O_D <= 32'b00111111011111100000000000000000;//1-2^(-5-2)
            5'b00010: O_D <= 32'b00111111011111000000000000000000;//1-2^(-4-2)   
            5'b00011: O_D <= 32'b00111111011110000000000000000000;//1-2^(-3-2) 
            5'b00100: O_D <= 32'b00111111011100000000000000000000;//1-2^(-2-2) 
            5'b00101: O_D <= 32'b00111111011000000000000000000000;//1-2^(-1-2) 
            5'b00110: O_D <= 32'b00111111010000000000000000000000;//1-2^(-0-2) 
            5'b00111: O_D <= 32'b00111111000000000000000000000000;//2^(-1) 
            5'b01000: O_D <= 32'b00111110100000000000000000000000;//2^(-2) 
            5'b01001: O_D <= 32'b00111110000000000000000000000000;//2^(-3) 
            5'b01010: O_D <= 32'b00111101100000000000000000000000;//2^(-4) 
            5'b01011: O_D <= 32'b00111101100000000000000000000000;//2^(-4) 
            5'b01100: O_D <= 32'b00111101000000000000000000000000;//2^(-5) 
            5'b01101: O_D <= 32'b00111100100000000000000000000000;//2^(-6) 
            5'b01110: O_D <= 32'b00111100000000000000000000000000;//2^(-7) 
            5'b01111: O_D <= 32'b00111100000000000000000000000000;//2^(-7) 
            5'b10000: O_D <= 32'b00111011100000000000000000000000;//2^(-8) 
            5'b10001: O_D <= 32'b00111011000000000000000000000000;//2^(-9) 
            5'b10010: O_D <= 32'b00111010100000000000000000000000;//2^(-10) 
            5'b10011: O_D <= 32'b00111010000000000000000000000000;//2^(-11) 
            5'b10100: O_D <= 32'b00111010000000000000000000000000;//2^(-11) 
            5'b10101: O_D <= 32'b00111001100000000000000000000000;//2^(-12) 
            5'b10110: O_D <= 32'b00111001000000000000000000000000;//2^(-13) 
            5'b10111: O_D <= 32'b00111000011111111111111111111110;//2^(-14) 
            5'b11000: O_D <= 32'b00111000011111111111111111111110;//2^(-14) 
            5'b11001: O_D <= 32'b00110111111111111111111111111100;//2^(-15) 
            5'b11010: O_D <= 32'b00110111011111111111111111110110;//2^(-16) 
            5'b11011: O_D <= 32'b00110111011111111111111111110110;//2^(-16) 
            5'b11100: O_D <= 32'b00110110111111111111111111110110;//2^(-17) 
            5'b11101: O_D <= 32'b00110110011111111111111111100000;//2^(-18) 
            5'b11110: O_D <= 32'b00110110011111111111111111100000;//2^(-18) 
            5'b11111: O_D <= 32'b00110101111111111111111110110100;//2^(-19) 
            default:  O_D <= 32'b00000000000000000000000000000000;
        endcase
        
endmodule