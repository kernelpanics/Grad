`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 06/29/2016 07:18:32 PM
// Design Name: 
// Module Name: Priority_Encoder
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module Priority_Encoder (

   input wire [31:0] d_in,
   output wire [7:0] d_out
   ); 

    assign d_out = (d_in[31]==1'b1) ? 8'b00011111:                  
                   (d_in[30]==1'b1) ? 8'b00011110:
                   (d_in[29]==1'b1) ? 8'b00011101:
                   (d_in[28]==1'b1) ? 8'b00011100:
                   (d_in[27]==1'b1) ? 8'b00011011:
                   (d_in[26]==1'b1) ? 8'b00011010:
                   (d_in[25]==1'b1) ? 8'b00011001:
                   (d_in[24]==1'b1) ? 8'b00011000:
                   (d_in[23]==1'b1) ? 8'b00010111:
                   (d_in[22]==1'b1) ? 8'b00010110:
                   (d_in[21]==1'b1) ? 8'b00010101:
                   (d_in[20]==1'b1) ? 8'b00010100:
                   (d_in[19]==1'b1) ? 8'b00010011:
                   (d_in[18]==1'b1) ? 8'b00010010:
                   (d_in[17]==1'b1) ? 8'b00010001:
                   (d_in[16]==1'b1) ? 8'b00010000:
                   (d_in[15]==1'b1) ? 8'b00001111:
                   (d_in[14]==1'b1) ? 8'b00001110:
                   (d_in[13]==1'b1) ? 8'b00001101:
                   (d_in[12]==1'b1) ? 8'b00001100:
                   (d_in[11]==1'b1) ? 8'b00001011:
                   (d_in[10]==1'b1) ? 8'b00001010:
                   (d_in[9]==1'b1)  ? 8'b00001001:
                   (d_in[8]==1'b1)  ? 8'b00001000: 
                   (d_in[7]==1'b1)  ? 8'b00000111:
                   (d_in[6]==1'b1)  ? 8'b00000110:
                   (d_in[5]==1'b1)  ? 8'b00000101:
                   (d_in[4]==1'b1)  ? 8'b00000100:
                   (d_in[3]==1'b1)  ? 8'b00000011:
                   (d_in[2]==1'b1)  ? 8'b00000010:
                   (d_in[1]==1'b1)  ? 8'b00000001: 8'b00000000;
                           
endmodule